library verilog;
use verilog.vl_types.all;
entity InterConn_Multiplexer is
    port(
        bus_grant       : in     vl_logic_vector(1 downto 0);
        slave_select    : in     vl_logic_vector(1 downto 0);
        M1_RX_DATA      : out    vl_logic;
        M1_SLAVE_VALID  : out    vl_logic;
        M1_SLAVE_READY  : out    vl_logic;
        M1_CLK          : in     vl_logic;
        M1_RST          : in     vl_logic;
        M1_VALID        : in     vl_logic;
        M1_TX_ADDR      : in     vl_logic;
        M1_TX_DATA      : in     vl_logic;
        M1_WRITE_EN     : in     vl_logic;
        M1_READ_EN      : in     vl_logic;
        M1_READY        : in     vl_logic;
        M1_TX_BURST     : in     vl_logic;
        M2_RX_DATA      : out    vl_logic;
        M2_SLAVE_VALID  : out    vl_logic;
        M2_SLAVE_READY  : out    vl_logic;
        M2_CLK          : in     vl_logic;
        M2_RST          : in     vl_logic;
        M2_VALID        : in     vl_logic;
        M2_TX_ADDR      : in     vl_logic;
        M2_TX_DATA      : in     vl_logic;
        M2_WRITE_EN     : in     vl_logic;
        M2_READ_EN      : in     vl_logic;
        M2_READY        : in     vl_logic;
        M2_TX_BURST     : in     vl_logic;
        S1_DATA_TX      : in     vl_logic;
        S1_SLAVE_READY  : in     vl_logic;
        S1_SLAVE_VALID  : in     vl_logic;
        S1_CLK          : out    vl_logic;
        S1_RST          : out    vl_logic;
        S1_M_VALID      : out    vl_logic;
        S1_M_READY      : out    vl_logic;
        S1_RX_ADDR      : out    vl_logic;
        S1_RX_DATA      : out    vl_logic;
        S1_WRITE_EN     : out    vl_logic;
        S1_READ_EN      : out    vl_logic;
        S1_RX_BURST     : out    vl_logic;
        S2_DATA_TX      : in     vl_logic;
        S2_SLAVE_READY  : in     vl_logic;
        S2_SLAVE_VALID  : in     vl_logic;
        S2_CLK          : out    vl_logic;
        S2_RST          : out    vl_logic;
        S2_M_VALID      : out    vl_logic;
        S2_M_READY      : out    vl_logic;
        S2_RX_ADDR      : out    vl_logic;
        S2_RX_DATA      : out    vl_logic;
        S2_WRITE_EN     : out    vl_logic;
        S2_READ_EN      : out    vl_logic;
        S2_RX_BURST     : out    vl_logic;
        S3_DATA_TX      : in     vl_logic;
        S3_SLAVE_READY  : in     vl_logic;
        S3_SLAVE_VALID  : in     vl_logic;
        S3_CLK          : out    vl_logic;
        S3_RST          : out    vl_logic;
        S3_M_VALID      : out    vl_logic;
        S3_M_READY      : out    vl_logic;
        S3_RX_ADDR      : out    vl_logic;
        S3_RX_DATA      : out    vl_logic;
        S3_WRITE_EN     : out    vl_logic;
        S3_READ_EN      : out    vl_logic;
        S3_RX_BURST     : out    vl_logic
    );
end InterConn_Multiplexer;
