

module input_commands #(parameter SLAVE_LEN=2, parameter ADDR_LEN=12, parameter DATA_LEN=8, parameter BURST_LEN=12)(
	input logic clk, 
	input logic reset,
	
	input logic button1,
	input logic button2,
	input logic button3,
	input logic [ADDR_LEN-1:0]switch_array,
	input logic mode_switch,
	input logic rw_switch1,
	input logic rw_switch2,


	output logic read1,
	output logic write1,
	output logic [DATA_LEN-1:0]data1 = 0,
	output logic [ADDR_LEN:0]address1 = 0,
	output logic [SLAVE_LEN-1:0]slave1 = 1,
	output logic [BURST_LEN:0]burst_num1 = 0,
	output logic read2,
	output logic write2,
	output logic [DATA_LEN-1:0]data2 = 0,
	output logic [ADDR_LEN:0]address2 = 0,
	output logic [SLAVE_LEN-1:0]slave2 = 1,
	output logic [BURST_LEN:0]burst_num2 = 0);
	
logic [2:0]config_state = 0;
logic [1:0]master = 1;
logic [DATA_LEN-1:0]data = 0;
logic [ADDR_LEN:0]address = 0;
logic [SLAVE_LEN-1:0]slave = 1;
logic [BURST_LEN:0]burst_num = 1;

logic button1_old = 0;
logic button2_old = 0;
logic button3_old = 0;
logic button1_edge;
logic button2_edge;
logic button3_edge;
assign button1_edge = (button1_old == 0 && button1 == 1) ? 1 : 0;
assign button2_edge = (button2_old == 0 && button2 == 1) ? 1 : 0;
assign button3_edge = (button3_old == 0 && button3 == 1) ? 1 : 0;

always @(posedge clk)
begin
	button1_old <= button1;
	button2_old <= button2;
	button3_old <= button3;
end

parameter SLAVE_NUM = 3;
parameter BURST_MAX = 12'hFFF;


parameter IDLE_CONFIG=0, SELECT_MASTER=1, SELECT_SLAVE=2, SELECT_ADDRESS=3, SELECT_DATA=4,
				SELECT_BURST=5, FINISH=6;
				
//wire [3:0]display_val1;
//wire [3:0]display_val2;
//wire [3:0]display_val3;
//wire [3:0]display_val4;

//assign display_val1 = (mode_switch == 0)?(
//							(config_state==1)?{2'b00,master}:
//							(config_state==2)?{2'b00,slave}:
//							(config_state==3)?switch_array[3:0]:
//							(config_state==4)?switch_array[3:0]:
//							(config_state==5)?switch_array[3:0]:0):0;
//							
//assign display_val2 = (mode_switch == 0)?(
//							(config_state==3)?switch_array[7:4]:
//							(config_state==4)?switch_array[7:4]:
//							(config_state==5)?switch_array[7:4]:0):0;
//							
//assign display_val3 = (mode_switch == 0)?(
//							(config_state==3)?switch_array[11:8]:
//							(config_state==5)?switch_array[11:8]:0):0;
//							
//assign display_val4 = (mode_switch == 0)?{1'b0,config_state}:0;
				
				
assign read1 = (mode_switch==1 && rw_switch1==1) ? button1 : 0;
assign write1 = (mode_switch==1 && rw_switch1==0) ? button1 : 0;

assign read2 = (mode_switch==1 && rw_switch2==1) ? button2 : 0;
assign write2 = (mode_switch==1 && rw_switch2==0) ? button2 : 0;


always @ (posedge reset or posedge clk)//button1 or posedge button2 or posedge button3 or posedge mode_switch) 
begin
	if (reset)
	begin
		config_state <= IDLE_CONFIG;
		master <= 1;
		slave <= 1;
		address <= 0;
		data <= 0;
		burst_num <= 1;
		slave1 <= 1;
		address1 <= 0;
		data1 <= 0;
		burst_num1 <= 1;
		slave2 <= 1;
		address2 <= 0;
		data2 <= 0;
		burst_num2 <= 1;
	end	
	
	else
	begin
		if (mode_switch==1)
		begin
			config_state <= IDLE_CONFIG;
			master <= 1;
			slave <= 1;
			address <= 0;
			data <= 0;
			burst_num <= 1;
		end
		else
		begin
		
			case(config_state)	
			
			IDLE_CONFIG:
			begin
				if (button1_edge==1 || button2_edge==1 || button3_edge==1)
				begin
					config_state <= SELECT_MASTER;
				end
				else
				begin
					config_state <= IDLE_CONFIG;
				end
				master <= 1;
				slave <= 1;
				address <= 0;
				data <= 0;
				burst_num <= 1;
				slave1 <= slave1;
				address1 <= address1;
				data1 <= data1;
				burst_num1 <= burst_num1;
				slave2 <= slave2;
				address2 <= address2;
				data2 <= data2;
				burst_num2 <= burst_num2;
			end
			
			SELECT_MASTER:
			begin
				if (button3_edge==1)     //button3 - KEY2
				begin
					config_state <= SELECT_SLAVE;
					master<=master;
				end
				else
				begin
					config_state <= SELECT_MASTER;
					if (button1_edge==1)    //button1 - KEY1 
					begin
						if (master==1)
							master <= 2;
						else
							master <= 1;
					end
					else if (button2_edge==1)  //button2 - KEY0
					begin
						if (master==1)
							master <= 2;
						else
							master <= 1;
					end
					else
					begin
						master<=master;
					end
				end
				slave <= slave;
				address <= address;
				data <= data;
				burst_num <= burst_num;
				slave1 <= slave1;
				address1 <= address1;
				data1 <= data1;
				burst_num1 <= burst_num1;
				slave2 <= slave2;
				address2 <= address2;
				data2 <= data2;
				burst_num2 <= burst_num2;
			end
			
			SELECT_SLAVE:
			begin
				if (button3_edge==1)
				begin
					config_state <= SELECT_ADDRESS;
					slave<=slave;
				end
				else
				begin
					config_state <= SELECT_SLAVE;
					if (button1_edge==1)
					begin
						if (slave>=SLAVE_NUM)
							slave <= 0;
						else
							slave <= slave+1;
					end
					else if (button2_edge==1)
					begin
						if (slave==1)
							slave <= SLAVE_NUM;
						else
							slave <= slave-1;
					end
					else
					begin
						slave<=slave;
					end
				end
				master <= master;
				address <= address;
				data <= data;
				burst_num <= burst_num;
				slave1 <= slave1;
				address1 <= address1;
				data1 <= data1;
				burst_num1 <= burst_num1;
				slave2 <= slave2;
				address2 <= address2;
				data2 <= data2;
				burst_num2 <= burst_num2;
			end
			
			SELECT_ADDRESS:
			begin
				if (button1_edge==1 || button2_edge==1 || button3_edge==1)
				begin
					config_state <= SELECT_DATA;
					address <= switch_array;
				end
				else
				begin
					config_state <= SELECT_ADDRESS;
					address <= address;
				end
				master <= master;
				slave <= slave;
				data <= data;
				burst_num <= burst_num;
				slave1 <= slave1;
				address1 <= address1;
				data1 <= data1;
				burst_num1 <= burst_num1;
				slave2 <= slave2;
				address2 <= address2;
				data2 <= data2;
				burst_num2 <= burst_num2;
			end
			
			SELECT_DATA:
			begin
				if (button1_edge==1 || button2_edge==1 || button3_edge==1)
				begin
					config_state <= SELECT_BURST;
					data <= switch_array[7:0];
				end
				else
				begin
					config_state <= SELECT_DATA;
					data <= data;
				end
				master <= master;
				slave <= slave;
				address <= address;
				burst_num <= burst_num;
				slave1 <= slave1;
				address1 <= address1;
				data1 <= data1;
				burst_num1 <= burst_num1;
				slave2 <= slave2;
				address2 <= address2;
				data2 <= data2;
				burst_num2 <= burst_num2;
			end
				
			SELECT_BURST:
			begin
				if (button1_edge==1 || button2_edge==1 || button3_edge==1)
				begin
					config_state <= FINISH;
					if (switch_array >= BURST_MAX)
						burst_num <= BURST_MAX;
					else
						burst_num <= switch_array;
				end
				else
				begin
					config_state <= SELECT_BURST;
					burst_num <= burst_num;
				end
				master <= master;
				slave <= slave;
				address <= address;
				data <= data;
				slave1 <= slave1;
				address1 <= address1;
				data1 <= data1;
				burst_num1 <= burst_num1;
				slave2 <= slave2;
				address2 <= address2;
				data2 <= data2;
				burst_num2 <= burst_num2;
			end
		
			FINISH:
			begin
				if (button1_edge==1 || button2_edge==1 || button3_edge==1)
				begin
					config_state <= IDLE_CONFIG;
					if (master==1)
					begin
						slave1 <= slave;
						address1 <= address;
						data1 <= data;
						burst_num1 <= burst_num;
						slave2 <= slave2;
						address2 <= address2;
						data2 <= data2;
						burst_num2 <= burst_num2;
					end
					else
					begin
						slave1 <= slave1;
						address1 <= address1;
						data1 <= data1;
						burst_num1 <= burst_num1;
						slave2 <= slave;
						address2 <= address;
						data2 <= data;
						burst_num2 <= burst_num;
					end
					master <= 1;
					slave <= 1;
					address <= 0;
					data <= 0;
					burst_num <= 1;
				end
				else
				begin
					config_state <= FINISH;
					master <= master;
					slave <= slave;
					address <= address;
					data <= data;
					burst_num <= burst_num;
					slave1 <= slave1;
					address1 <= address1;
					data1 <= data1;
					burst_num1 <= burst_num1;
					slave2 <= slave2;
					address2 <= address2;
					data2 <= data2;
					burst_num2 <= burst_num2;
				end
			end
		
			default:
			begin
				config_state <= IDLE_CONFIG;
				master <= 1;
				slave <= 1;
				address <= 0;
				data <= 0;
				burst_num <= 1;
				slave1 <= 1;
				address1 <= 0;
				data1 <= 0;
				burst_num1 <= 1;
				slave2 <= 1;
				address2 <= 0;
				data2 <= 0;
				burst_num2 <= 1;
			end
			endcase
		end
		
	end
end


endmodule