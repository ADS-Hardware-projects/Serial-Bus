//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Saliya Dinusha
// 
// Create Date: 10/06/2023 03:36:17 PM
// Design Name: 
// Module Name: master_in_port_tb
// Project Name: SystemBus
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: NO
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module master_in_port#(parameter WORD_SIZE=8, parameter BURST_SIZE=15 )(

    //global inputs
    input logic clk,
    input logic rst,

    //inputs from bus side
    input logic rx_data,
    input logic s_valid,
	 input logic tx_done,

    //inputs from master core side
    input logic [1:0] instruction,
    input logic [BURST_SIZE-1:0] burst_size,

	 //outputs to bus side
    output logic m_ready,

    
    //outputs to master core side
    output logic rx_done,
    output logic [WORD_SIZE-1:0] s_data,
    output logic new_data


);

    logic [2:0] state= 3'b000;
    logic [WORD_SIZE-1:0] temp_data;
    parameter IDLE=0, READ= 1, RECIEVE = 2;

    integer bit_count =0;
    integer burst_count = 0;

    always @ (posedge clk or posedge rst) 
    begin

        if (rst)
        begin
            bit_count<=0;
            burst_count<=0;
            s_data <=0;
            temp_data<= 0;
            m_ready <= 1;
            state <= IDLE;
            rx_done <= 0;
				new_data <= 0;
        end
        else
        begin
            case (state)

            IDLE:
            begin
                if (instruction== 2'b11 && tx_done == 1)
                begin
							bit_count<=0;
							burst_count<=0;
							s_data <= s_data;
							temp_data<= temp_data;
							m_ready <= 1;
							state <= READ;
							rx_done <= 0;
							new_data <= 0;

                end
                else
                begin
							bit_count<= bit_count;
							burst_count<= burst_count;
							s_data <= s_data;
							temp_data<= temp_data;
							m_ready <= 1;
							state <= IDLE;
							rx_done <= 0;
							new_data <= 0;
                end
            end

            READ:
            begin
                if (m_ready==1 && s_valid == 1)
                begin
                    state <= RECIEVE;
                    m_ready <= 0;
                    new_data <=0;

                end
                else
                begin
                    state = READ;
                end

            end


            RECIEVE:
            begin

                if (bit_count >= WORD_SIZE-1)
                begin

                    bit_count <= 0;
                    new_data <= 1;
                    temp_data[bit_count] <= rx_data;
                    
                    m_ready <= 1;
                    s_data[bit_count] <= rx_data;
                    s_data[WORD_SIZE-2:0]<= temp_data[WORD_SIZE-2:0];

                    if (burst_count>= burst_size-1)
                    begin
                        state <= IDLE;
                        rx_done <= 1;
                        burst_count <=0;
                        
                    end

                    else
                    begin
                        burst_count <= burst_count+1;
                        state <= RECIEVE;
                        m_ready <= 0;
                        rx_done <= 0;
                        
                    end

                end

                else
                begin
                    temp_data[bit_count] <= rx_data;
                    bit_count <= bit_count + 1;
                    state <= RECIEVE;
                    new_data <= 0;

                end

            end
            endcase
        end

    end


endmodule